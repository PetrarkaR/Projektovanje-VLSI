LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE DEFS IS
	CONSTANT load : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("00000");
	CONSTANT setf : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("00001");
	CONSTANT clrf : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("00010");
	CONSTANT add : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("00011");
	CONSTANT addc : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("00100");
	CONSTANT sub_op : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("00101");
	CONSTANT subc : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("00110");
	CONSTANT rol_op : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("00111");
	CONSTANT rolc : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("01000");
	CONSTANT ror_op : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("01001");
	CONSTANT rorc : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("01010");
	CONSTANT and_op : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("01011");
	CONSTANT or_op : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("01100");
	CONSTANT xor_op : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("01101");
	CONSTANT not_op : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("01110");
	CONSTANT loadl : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("01111");
	CONSTANT store : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("10000");
	CONSTANT read : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("10001");
	CONSTANT write : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("10010");
	CONSTANT jnf : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("10011");
	CONSTANT jf : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("10100");
	CONSTANT jnz : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("10101");
	CONSTANT jz : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("10110");
	CONSTANT jmp : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("10111");
	CONSTANT nop : STD_LOGIC_VECTOR(4 DOWNTO 0) := ("11000");
END PACKAGE DEFS;